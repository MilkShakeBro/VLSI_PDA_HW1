/users/student/mr112/whhung23/HW1/NangateOpenCellLibrary.lef